** sch_path: /foss/designs/eda/designs/gmid/vt_W_n.sch
**.subckt vt_W_n
Xm1 d g GND b sg13_lv_nmos W={Wx} L={Lx} ng={nx} m=1
Vgs g GND 0.6
Vds d GND 0.6
Vsb GND b {vsbx}
**** begin user architecture code
 .lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt



.param temp=27
.param Wx=5u
.param Lx=0.13u
.param nx=1
.param Vsbx=0
.dc Vds 0.6 1.2 0.6
.save @n.xm1.nsg13_lv_nmos[vth]
.save @n.xm1.nsg13_lv_nmos[ids]


.control
*pre_osdi ./psp103_nqs.osdi
set wr_singlescale
*set wr_vecnames
option numdgt = 3

foreach W_val 0.15u 0.25u 0.35u 0.45u 0.55u 0.65u 0.75u 0.85u 0.95u
+ 1u 2u 3u 4u 5u 6u 7u 8u 9u 10u 11u 12u 13u 14u 15u 16u 17u 18u 19u 20u
+ 25u 30u 35u 40u 45u 50u
  alterparam Wx = $W_val
  reset
  run
  wrdata vt_W_n.txt all
  destroy $curplot
  set appendwrite
end
* show
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
